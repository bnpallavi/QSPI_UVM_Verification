class qspi_sequencer extends uvm_sequencer #(qspi_item);

   `uvm_component_utils(qspi_sequencer)

   function new(string name, uvm_component parent);
      super.new(name,parent);
   endfunction

endclass
